* SPICE3 file created from CVBT.ext - technology: scmos

.option scale=0.3u

