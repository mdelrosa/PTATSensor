magic
tech scmos
timestamp 1415294909
<< nwell >>
rect 9 9 47 47
<< pdiffusion >>
rect 22 33 34 34
rect 22 23 23 33
rect 33 23 34 33
rect 22 22 34 23
<< pdcontact >>
rect 23 23 33 33
<< psubstratepdiff >>
rect 0 55 56 56
rect 0 51 1 55
rect 55 51 56 55
rect 0 50 56 51
rect 0 48 6 50
rect 0 8 1 48
rect 5 8 6 48
rect 50 48 56 50
rect 50 37 51 48
rect 55 37 56 48
rect 50 20 56 37
rect 0 6 6 8
rect 50 8 51 20
rect 55 8 56 20
rect 50 6 56 8
rect 0 5 56 6
rect 0 1 1 5
rect 55 1 56 5
rect 0 0 56 1
<< nsubstratendiff >>
rect 12 43 44 44
rect 12 39 13 43
rect 43 39 44 43
rect 12 38 44 39
rect 12 36 18 38
rect 12 20 13 36
rect 17 20 18 36
rect 38 36 44 38
rect 38 30 39 36
rect 43 30 44 36
rect 12 18 18 20
rect 38 18 44 30
rect 12 17 44 18
rect 12 13 13 17
rect 43 13 44 17
rect 12 12 44 13
<< psubstratepcontact >>
rect 1 51 55 55
rect 1 8 5 48
rect 51 37 55 48
rect 51 8 55 20
rect 1 1 55 5
<< nsubstratencontact >>
rect 13 39 43 43
rect 13 20 17 36
rect 39 30 43 36
rect 13 13 43 17
<< metal1 >>
rect 1 48 5 51
rect 51 48 55 51
rect 13 36 17 39
rect 39 36 43 39
rect 55 37 59 41
rect 43 30 59 34
rect 33 23 59 27
rect 13 17 17 20
rect 1 5 5 8
rect 51 5 55 8
<< labels >>
rlabel metal1 58 38 59 40 3 C
rlabel metal1 58 31 59 33 3 B
rlabel metal1 58 24 59 26 3 E
<< end >>
