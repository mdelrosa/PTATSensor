magic
tech scmos
timestamp 1411404921
<< ntransistor >>
rect 8 7 10 11
<< ptransistor >>
rect 8 23 10 27
<< ndiffusion >>
rect 7 7 8 11
rect 10 7 11 11
<< pdiffusion >>
rect 7 23 8 27
rect 10 23 11 27
<< ndcontact >>
rect 3 7 7 11
rect 11 7 15 11
<< pdcontact >>
rect 3 23 7 27
rect 11 23 15 27
<< polysilicon >>
rect 8 27 10 29
rect 8 11 10 23
rect 8 5 10 7
<< polycontact >>
rect 4 15 8 19
<< metal1 >>
rect 3 27 7 31
rect 11 19 15 23
rect 0 15 4 19
rect 11 15 18 19
rect 11 11 15 15
rect 3 3 7 7
<< m2contact >>
rect 3 31 7 35
rect 3 -1 7 3
<< metal2 >>
rect 0 38 3 43
rect 0 35 18 38
rect 0 31 3 35
rect 7 31 18 35
rect 0 -1 3 3
rect 7 -1 18 3
rect 0 -4 18 -1
rect 0 -5 3 -4
<< labels >>
rlabel metal1 15 15 18 19 7 out
rlabel metal2 0 31 18 35 5 Vdd
rlabel metal2 0 -1 18 3 1 GND
rlabel metal1 0 15 4 19 3 in
<< end >>
