magic
tech scmos
timestamp 1418517441
<< ntransistor >>
rect -6 -105 394 -101
rect 399 -105 429 -101
rect -45 -513 -41 -113
rect -1 -512 3 -113
rect 311 -244 411 -234
<< ptransistor >>
rect 108 -46 138 -36
rect 156 -46 166 -36
rect 175 -46 185 -36
rect 191 -46 204 -36
<< ndiffusion >>
rect -6 -96 394 -95
rect -6 -100 -5 -96
rect 393 -100 394 -96
rect -6 -101 394 -100
rect 399 -96 429 -95
rect 399 -100 401 -96
rect 427 -100 429 -96
rect 399 -101 429 -100
rect -49 -102 -37 -101
rect -49 -110 -48 -102
rect -38 -110 -37 -102
rect -49 -111 -37 -110
rect -45 -113 -41 -111
rect -6 -106 394 -105
rect -6 -110 -5 -106
rect 393 -110 394 -106
rect -6 -111 394 -110
rect 399 -106 429 -105
rect 399 -110 401 -106
rect 427 -110 429 -106
rect 399 -111 429 -110
rect -1 -113 3 -111
rect 311 -225 411 -223
rect 311 -233 313 -225
rect 409 -233 411 -225
rect 311 -234 411 -233
rect 311 -246 411 -244
rect 311 -254 313 -246
rect 409 -254 411 -246
rect 311 -255 411 -254
rect -45 -515 -41 -513
rect -1 -514 3 -512
rect -5 -515 7 -514
rect -49 -516 -37 -515
rect -49 -520 -48 -516
rect -38 -520 -37 -516
rect -5 -519 -4 -515
rect 6 -519 7 -515
rect -5 -520 7 -519
rect -49 -521 -37 -520
<< pdiffusion >>
rect 156 -30 166 -29
rect 108 -31 138 -30
rect 108 -35 109 -31
rect 137 -35 138 -31
rect 108 -36 138 -35
rect 156 -35 157 -30
rect 165 -35 166 -30
rect 156 -36 166 -35
rect 175 -30 185 -29
rect 175 -35 176 -30
rect 184 -35 185 -30
rect 175 -36 185 -35
rect 191 -30 204 -29
rect 191 -35 192 -30
rect 203 -35 204 -30
rect 191 -36 204 -35
rect 108 -47 138 -46
rect 108 -51 109 -47
rect 137 -51 138 -47
rect 108 -52 138 -51
rect 156 -48 166 -46
rect 156 -53 157 -48
rect 165 -53 166 -48
rect 156 -54 166 -53
rect 175 -48 185 -46
rect 175 -53 176 -48
rect 184 -53 185 -48
rect 175 -54 185 -53
rect 191 -48 204 -46
rect 191 -53 192 -48
rect 203 -53 204 -48
rect 191 -54 204 -53
<< ndcontact >>
rect -5 -100 393 -96
rect 401 -100 427 -96
rect -48 -110 -38 -102
rect -5 -110 393 -106
rect 401 -110 427 -106
rect 313 -233 409 -225
rect 313 -254 409 -246
rect -48 -520 -38 -516
rect -4 -519 6 -515
<< pdcontact >>
rect 109 -35 137 -31
rect 157 -35 165 -30
rect 176 -35 184 -30
rect 192 -35 203 -30
rect 109 -51 137 -47
rect 157 -53 165 -48
rect 176 -53 184 -48
rect 192 -53 203 -48
<< polysilicon >>
rect 105 -46 108 -36
rect 138 -46 156 -36
rect 166 -46 175 -36
rect 185 -46 191 -36
rect 204 -46 210 -36
rect 143 -48 151 -46
rect 143 -53 144 -48
rect 150 -53 151 -48
rect 143 -54 151 -53
rect 431 -95 438 -94
rect 431 -100 432 -95
rect 437 -100 438 -95
rect 431 -101 438 -100
rect -36 -103 -27 -102
rect -36 -109 -35 -103
rect -28 -109 -27 -103
rect -9 -105 -6 -101
rect 394 -105 399 -101
rect 429 -105 438 -101
rect -36 -113 -27 -109
rect -49 -513 -45 -113
rect -41 -512 -1 -113
rect 3 -234 7 -113
rect 3 -244 311 -234
rect 411 -244 414 -234
rect 3 -512 7 -244
rect -41 -513 -3 -512
<< polycontact >>
rect 144 -53 150 -48
rect 432 -100 437 -95
rect -35 -109 -28 -103
<< metal1 >>
rect 100 -31 157 -30
rect 100 -35 109 -31
rect 137 -35 157 -31
rect 165 -35 176 -30
rect 184 -35 192 -30
rect 203 -35 213 -30
rect -49 -51 109 -48
rect 176 -48 184 -47
rect 137 -51 138 -48
rect -49 -52 138 -51
rect -49 -102 -38 -52
rect 143 -53 144 -48
rect 150 -53 157 -48
rect 165 -53 166 -48
rect 156 -92 166 -53
rect 176 -73 184 -53
rect 191 -53 192 -48
rect 203 -53 454 -48
rect 191 -56 454 -53
rect 176 -83 427 -73
rect -5 -96 393 -92
rect 401 -95 427 -83
rect 401 -96 432 -95
rect 427 -100 432 -96
rect -5 -101 393 -100
rect -50 -110 -48 -102
rect -38 -103 -27 -102
rect -38 -109 -35 -103
rect -28 -109 -27 -103
rect -38 -110 -27 -109
rect -50 -111 -27 -110
rect 313 -225 460 -223
rect 409 -233 460 -225
rect 312 -254 313 -246
rect 312 -263 408 -254
rect 347 -515 372 -263
rect -49 -516 -29 -515
rect -49 -520 -48 -516
rect -38 -520 -29 -516
rect -18 -519 -4 -515
rect 6 -519 266 -515
rect -18 -520 266 -519
rect 277 -520 372 -515
rect 347 -523 372 -520
<< m2contact >>
rect 93 -35 100 -30
rect 213 -35 220 -30
rect -29 -523 -18 -515
rect 266 -523 277 -515
<< metal2 >>
rect -59 -30 454 -27
rect -59 -35 93 -30
rect 100 -35 213 -30
rect 220 -35 454 -30
rect -59 -36 454 -35
rect -50 -515 483 -514
rect -50 -523 -29 -515
rect -18 -523 266 -515
rect 277 -523 483 -515
rect -50 -524 483 -523
<< labels >>
rlabel metal1 455 -231 458 -224 1 I_pull
rlabel metal2 449 -35 452 -28 5 Vdd
rlabel metal1 449 -55 452 -49 1 I_push
rlabel metal2 478 -522 481 -515 7 Gnd
<< end >>
