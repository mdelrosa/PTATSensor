magic
tech scmos
timestamp 1418693430
<< electrodecontact >>
rect 78 792 86 800
rect 115 792 123 800
rect 176 792 184 800
rect 216 792 224 800
rect 278 792 286 800
rect 317 792 325 800
rect 378 792 386 800
rect 417 792 425 800
rect 480 792 488 800
rect 520 792 528 800
rect 582 792 590 800
rect 620 792 628 800
rect 78 753 86 761
rect 78 692 85 699
rect 115 692 122 699
rect 176 692 184 700
rect 217 692 225 700
rect 277 692 285 700
rect 317 692 325 700
rect 378 692 386 700
rect 417 692 425 700
rect 480 692 488 700
rect 519 692 527 700
rect 583 692 591 700
rect 620 692 628 700
rect 78 656 85 663
rect 482 657 490 665
rect 520 657 528 665
rect 583 657 591 665
rect 620 657 628 665
rect 13 598 22 606
rect 78 595 85 602
rect 120 595 127 602
rect 178 595 185 602
rect 223 595 230 602
rect 381 595 388 602
rect 422 557 429 564
rect 482 557 489 564
rect 519 557 526 564
rect 583 557 590 564
rect 621 557 628 564
rect 423 537 429 543
rect 17 513 23 519
rect 78 496 85 503
rect 121 496 128 503
rect 179 496 186 503
rect 219 496 226 503
rect 280 496 287 503
rect 321 457 328 464
rect 484 454 491 461
rect 521 454 528 461
rect 584 454 591 461
rect 619 454 626 461
rect 80 390 87 397
rect 114 390 121 397
rect 181 390 188 397
rect 215 390 222 397
rect 619 392 626 398
rect 80 357 87 364
rect 584 357 591 364
rect 619 357 626 364
rect 79 290 86 297
rect 115 290 122 297
rect 181 290 188 297
rect 215 290 222 297
rect 281 290 288 297
rect 316 290 323 297
rect 382 291 389 298
rect 419 291 426 298
rect 484 291 491 298
rect 519 291 526 298
rect 584 291 591 298
rect 619 291 626 298
rect 79 256 86 263
rect 114 256 121 263
rect 181 256 188 263
rect 215 256 222 263
rect 281 255 288 262
rect 317 255 324 262
rect 382 255 389 262
rect 419 255 426 262
rect 484 255 491 262
rect 519 255 526 262
rect 583 255 590 262
rect 619 255 626 262
rect 13 192 19 198
<< electrodecap >>
rect 11 787 89 865
rect 112 787 190 865
rect 213 787 291 865
rect 314 787 392 865
rect 415 787 493 865
rect 516 787 594 865
rect 617 787 695 865
rect 11 688 89 766
rect 112 688 190 766
rect 213 688 291 766
rect 314 688 392 766
rect 415 688 493 766
rect 516 688 594 766
rect 617 688 695 766
rect 11 589 89 667
rect 112 589 190 667
rect 213 589 291 667
rect 314 589 392 667
rect 415 589 493 667
rect 516 589 594 667
rect 617 589 695 667
rect 11 489 89 567
rect 112 489 190 567
rect 213 489 291 567
rect 415 489 493 567
rect 516 489 594 567
rect 617 489 695 567
rect 11 388 89 466
rect 112 388 190 466
rect 213 388 291 466
rect 314 388 392 466
rect 415 388 493 466
rect 516 388 594 466
rect 617 388 695 466
rect 11 288 89 366
rect 112 288 190 366
rect 213 288 291 366
rect 314 288 392 366
rect 415 288 493 366
rect 516 288 594 366
rect 617 288 695 366
rect 11 187 89 265
rect 112 187 190 265
rect 213 187 291 265
rect 314 187 392 265
rect 415 187 493 265
rect 516 187 594 265
rect 617 187 695 265
<< ntransistor >>
rect -85 110 -79 116
rect -65 110 -59 116
rect -80 52 -74 58
rect -19 52 -13 58
rect -89 21 -83 27
rect -28 21 -22 27
<< ndiffusion >>
rect -85 116 -79 118
rect -65 116 -59 118
rect -85 107 -79 110
rect -65 107 -59 110
rect -81 52 -80 58
rect -74 52 -73 58
rect -20 52 -19 58
rect -13 52 -12 58
rect -99 21 -89 27
rect -83 21 -82 27
rect -32 21 -28 27
rect -22 21 -21 27
<< ndcontact >>
rect -85 118 -79 124
rect -65 118 -59 124
rect -85 101 -79 107
rect -65 101 -59 107
rect -87 52 -81 58
rect -73 52 -67 58
rect -26 52 -20 58
rect -12 52 -6 58
rect -105 21 -99 27
rect -82 21 -76 27
rect -38 21 -32 27
rect -21 21 -15 27
<< polysilicon >>
rect 4 865 702 872
rect 4 780 96 865
rect 105 780 197 865
rect 206 780 298 865
rect 307 780 399 865
rect 408 780 500 865
rect 509 780 601 865
rect 610 780 702 865
rect 610 773 617 780
rect 4 766 702 773
rect 4 681 96 766
rect 105 681 197 766
rect 206 681 298 766
rect 307 681 399 766
rect 408 681 500 766
rect 509 681 601 766
rect 610 681 702 766
rect 89 674 96 681
rect 610 674 617 681
rect 4 667 298 674
rect 4 588 96 667
rect 8 582 96 588
rect 105 582 197 667
rect 206 582 298 667
rect 307 589 399 674
rect 408 667 702 674
rect 307 582 394 589
rect 408 582 500 667
rect 509 582 601 667
rect 610 582 702 667
rect 4 531 96 574
rect 7 525 96 531
rect 4 489 96 525
rect 105 489 197 574
rect 206 489 298 574
rect 415 570 702 574
rect 408 566 702 570
rect 408 554 500 566
rect 411 548 500 554
rect 4 482 293 489
rect 408 482 500 548
rect 509 482 601 566
rect 610 555 702 566
rect 610 548 698 555
rect 610 482 702 548
rect 4 388 96 473
rect 105 388 197 473
rect 206 393 298 473
rect 314 468 399 473
rect 307 440 399 468
rect 307 433 395 440
rect 206 388 297 393
rect 4 381 297 388
rect 307 381 399 433
rect 408 388 500 473
rect 509 388 601 473
rect 610 388 702 473
rect 408 381 702 388
rect 4 373 11 381
rect 610 373 617 381
rect 4 288 96 373
rect 105 288 197 373
rect 206 288 298 373
rect 307 288 399 373
rect 408 288 500 373
rect 509 288 601 373
rect 610 288 702 373
rect 4 281 702 288
rect 610 272 617 281
rect 4 187 96 272
rect 105 187 197 272
rect 206 187 298 272
rect 307 187 399 272
rect 408 187 500 272
rect 509 187 601 272
rect 610 187 702 272
rect 4 186 702 187
rect 9 180 702 186
rect -299 121 -281 127
rect -150 121 -119 127
rect -170 110 -85 116
rect -79 110 -65 116
rect -59 110 -56 116
rect -298 76 -280 82
rect -151 76 -130 82
rect -80 58 -74 61
rect -19 58 -13 61
rect -80 47 -74 52
rect -19 47 -13 52
rect -89 27 -83 30
rect -28 27 -22 30
rect -89 18 -83 21
rect -28 18 -22 21
<< polycontact >>
rect 2 582 8 588
rect 394 582 401 589
rect 1 525 7 531
rect 408 570 415 577
rect 405 548 411 554
rect 293 482 300 489
rect 698 548 705 555
rect 307 468 314 475
rect 395 433 402 440
rect 3 180 9 186
rect -305 121 -299 127
rect -119 121 -113 127
rect -176 110 -170 116
rect -304 76 -298 82
rect -130 76 -124 82
rect -80 61 -74 67
rect -19 61 -13 67
rect -89 30 -83 36
rect -89 12 -83 18
rect -28 12 -22 18
<< metal1 >>
rect 86 792 115 800
rect 184 792 216 800
rect 286 792 317 800
rect 386 792 417 800
rect 488 792 520 800
rect 590 792 620 800
rect 78 761 86 792
rect 85 692 115 699
rect 184 692 217 700
rect 285 692 317 700
rect 386 692 417 700
rect 488 692 519 700
rect 591 692 620 700
rect 78 663 85 692
rect 620 665 628 692
rect 490 657 520 665
rect 591 657 620 665
rect -293 605 13 606
rect -286 598 13 605
rect 85 595 120 602
rect 185 595 223 602
rect 388 595 429 602
rect -39 582 2 588
rect 401 582 415 589
rect 408 577 415 582
rect 422 564 429 595
rect 489 557 519 564
rect 590 557 621 564
rect -79 548 405 554
rect 705 548 718 555
rect -70 537 423 543
rect -59 525 1 531
rect -48 513 17 519
rect 85 496 121 503
rect 186 496 219 503
rect 287 496 328 503
rect 300 482 314 489
rect 307 475 314 482
rect 321 464 328 496
rect 491 454 521 461
rect 591 454 619 461
rect 402 433 706 440
rect 87 390 114 397
rect 188 390 215 397
rect 80 364 87 390
rect 619 364 626 392
rect 591 357 619 364
rect 86 290 115 297
rect 188 290 215 297
rect 288 290 316 297
rect 389 291 419 298
rect 491 291 519 298
rect 591 291 619 298
rect 86 256 114 263
rect 188 256 215 263
rect 619 262 626 291
rect 288 255 317 262
rect 389 255 419 262
rect 491 255 519 262
rect 590 255 619 262
rect -139 192 13 198
rect -27 180 3 186
rect 725 168 1361 175
rect 713 154 1351 161
rect -106 140 -45 146
rect -113 121 -105 127
rect -305 110 -253 116
rect -177 110 -176 116
rect -286 69 -280 74
rect -151 69 -145 74
rect -130 18 -124 76
rect -112 67 -105 121
rect -85 124 -79 125
rect -65 124 -59 125
rect -79 101 -76 107
rect -59 101 -54 107
rect -85 98 -79 101
rect -85 92 -64 98
rect -94 82 -34 89
rect 1349 88 1361 95
rect -83 70 -13 76
rect -19 67 -13 70
rect -112 61 -80 67
rect -74 61 -73 67
rect 1349 58 1351 65
rect -95 52 -87 58
rect -27 52 -26 58
rect -73 49 -67 52
rect -12 49 -6 52
rect -73 43 -54 49
rect -48 44 6 49
rect -48 43 4 44
rect 0 41 4 43
rect -89 36 -83 37
rect -73 31 -64 37
rect -58 31 7 37
rect -73 27 -67 31
rect -21 27 -15 31
rect -106 21 -105 27
rect -76 21 -67 27
rect -39 21 -38 27
rect -130 12 -89 18
rect -67 12 -28 18
rect -81 0 1 7
<< m2contact >>
rect -293 598 -286 605
rect -45 582 -39 588
rect -85 548 -79 554
rect 718 548 725 555
rect -76 537 -70 543
rect -65 525 -59 531
rect -54 513 -48 519
rect 706 433 713 440
rect -145 192 -139 198
rect -33 180 -27 186
rect 718 168 725 175
rect 1361 168 1368 175
rect 706 154 713 161
rect 1351 154 1358 161
rect -112 140 -106 146
rect -45 140 -39 146
rect -253 110 -247 116
rect -183 110 -177 116
rect -292 69 -286 75
rect -145 69 -139 75
rect -85 125 -79 131
rect -65 125 -59 131
rect -76 101 -70 107
rect -54 101 -48 107
rect -64 92 -58 98
rect -101 82 -94 89
rect -34 82 -27 89
rect 1361 88 1368 95
rect -89 70 -83 76
rect -73 61 -67 67
rect 1351 58 1358 65
rect -101 52 -95 58
rect -33 52 -27 58
rect -54 43 -48 49
rect -89 37 -83 43
rect -64 31 -58 37
rect -112 21 -106 27
rect -45 21 -39 27
rect -73 12 -67 18
rect -88 0 -81 7
<< metal2 >>
rect -293 342 -286 598
rect -292 75 -286 342
rect -247 110 -183 116
rect -145 75 -139 192
rect -112 27 -106 140
rect -85 131 -79 548
rect -76 107 -70 537
rect -65 131 -59 525
rect -54 107 -48 513
rect -101 58 -95 82
rect -89 43 -83 70
rect -73 18 -67 61
rect -64 37 -58 92
rect -54 49 -48 101
rect -45 146 -39 582
rect -45 27 -39 140
rect -33 89 -27 180
rect 706 161 713 433
rect 718 175 725 548
rect -33 58 -27 82
rect 1351 65 1358 154
rect 1361 95 1368 168
rect -296 0 -268 5
rect -152 0 -88 5
use PTAT  PTAT_0
timestamp 1417640631
transform 1 0 -196 0 1 112
box -86 -112 61 38
use CMFFDiffAmp  CMFFDiffAmp_0
timestamp 1418250215
transform 1 0 661 0 1 50
box -661 -50 689 93
<< end >>
