magic
tech scmos
timestamp 1417680066
<< ptransistor >>
rect -17 -1 -11 5
rect -1 -1 5 5
rect 9 -1 15 5
rect 25 -1 31 5
rect 35 -1 41 5
rect 51 -1 57 5
rect 61 -1 67 5
rect 78 -1 84 5
rect 88 -1 94 5
rect 9 -24 15 -18
rect 35 -24 41 -18
rect 61 -24 67 -18
rect 88 -24 94 -18
rect 105 -24 111 -18
rect 115 -24 121 -18
<< pdiffusion >>
rect -17 11 -11 12
rect -17 7 -16 11
rect -12 7 -11 11
rect -17 5 -11 7
rect -1 11 5 12
rect -1 7 0 11
rect 4 7 5 11
rect -1 5 5 7
rect 9 11 15 12
rect 9 7 10 11
rect 14 7 15 11
rect 9 5 15 7
rect 25 11 31 12
rect 25 7 26 11
rect 30 7 31 11
rect 25 5 31 7
rect 35 11 41 12
rect 35 7 36 11
rect 40 7 41 11
rect 35 5 41 7
rect 51 11 57 12
rect 51 7 52 11
rect 56 7 57 11
rect 51 5 57 7
rect 61 11 67 12
rect 61 7 62 11
rect 66 7 67 11
rect 61 5 67 7
rect 78 11 84 12
rect 78 7 79 11
rect 83 7 84 11
rect 78 5 84 7
rect 88 11 94 12
rect 88 7 89 11
rect 93 7 94 11
rect 88 5 94 7
rect -17 -3 -11 -1
rect -17 -7 -16 -3
rect -12 -7 -11 -3
rect -17 -8 -11 -7
rect -1 -3 5 -1
rect -1 -7 0 -3
rect 4 -7 5 -3
rect -1 -8 5 -7
rect 9 -3 15 -1
rect 9 -7 10 -3
rect 14 -7 15 -3
rect 9 -8 15 -7
rect 25 -3 31 -1
rect 25 -7 26 -3
rect 30 -7 31 -3
rect 25 -8 31 -7
rect 35 -3 41 -1
rect 35 -7 36 -3
rect 40 -7 41 -3
rect 35 -8 41 -7
rect 51 -3 57 -1
rect 51 -7 52 -3
rect 56 -7 57 -3
rect 51 -8 57 -7
rect 61 -3 67 -1
rect 61 -7 62 -3
rect 66 -7 67 -3
rect 61 -8 67 -7
rect 78 -3 84 -1
rect 78 -7 79 -3
rect 83 -7 84 -3
rect 78 -8 84 -7
rect 88 -3 94 -1
rect 88 -7 89 -3
rect 93 -7 94 -3
rect 88 -8 94 -7
rect 9 -12 15 -11
rect 9 -16 10 -12
rect 14 -16 15 -12
rect 9 -18 15 -16
rect 35 -12 41 -11
rect 35 -16 36 -12
rect 40 -16 41 -12
rect 35 -18 41 -16
rect 61 -12 67 -11
rect 61 -16 62 -12
rect 66 -16 67 -12
rect 61 -18 67 -16
rect 88 -12 94 -11
rect 88 -16 89 -12
rect 93 -16 94 -12
rect 88 -18 94 -16
rect 105 -12 111 -11
rect 105 -16 106 -12
rect 110 -16 111 -12
rect 105 -18 111 -16
rect 115 -12 121 -11
rect 115 -16 116 -12
rect 120 -16 121 -12
rect 115 -18 121 -16
rect 9 -26 15 -24
rect 9 -30 10 -26
rect 14 -30 15 -26
rect 9 -31 15 -30
rect 35 -26 41 -24
rect 35 -30 36 -26
rect 40 -30 41 -26
rect 35 -31 41 -30
rect 61 -26 67 -24
rect 61 -30 62 -26
rect 66 -30 67 -26
rect 61 -31 67 -30
rect 88 -26 94 -24
rect 88 -30 89 -26
rect 93 -30 94 -26
rect 88 -31 94 -30
rect 105 -26 111 -24
rect 105 -30 106 -26
rect 110 -30 111 -26
rect 105 -31 111 -30
rect 115 -26 121 -24
rect 115 -30 116 -26
rect 120 -30 121 -26
rect 115 -31 121 -30
<< pdcontact >>
rect -16 7 -12 11
rect 0 7 4 11
rect 10 7 14 11
rect 26 7 30 11
rect 36 7 40 11
rect 52 7 56 11
rect 62 7 66 11
rect 79 7 83 11
rect 89 7 93 11
rect -16 -7 -12 -3
rect 0 -7 4 -3
rect 10 -7 14 -3
rect 26 -7 30 -3
rect 36 -7 40 -3
rect 52 -7 56 -3
rect 62 -7 66 -3
rect 79 -7 83 -3
rect 89 -7 93 -3
rect 10 -16 14 -12
rect 36 -16 40 -12
rect 62 -16 66 -12
rect 89 -16 93 -12
rect 106 -16 110 -12
rect 116 -16 120 -12
rect 10 -30 14 -26
rect 36 -30 40 -26
rect 62 -30 66 -26
rect 89 -30 93 -26
rect 106 -30 110 -26
rect 116 -30 120 -26
<< polysilicon >>
rect -28 4 -17 5
rect -28 0 -24 4
rect -20 0 -17 4
rect -28 -1 -17 0
rect -11 -1 -1 5
rect 5 -1 9 5
rect 15 -1 25 5
rect 31 -1 35 5
rect 41 -1 51 5
rect 57 -1 61 5
rect 67 -1 78 5
rect 84 -1 88 5
rect 94 -1 96 5
rect 7 -24 9 -18
rect 15 -24 35 -18
rect 41 -24 61 -18
rect 67 -24 88 -18
rect 94 -24 105 -18
rect 111 -24 115 -18
rect 121 -24 123 -18
<< polycontact >>
rect -24 0 -20 4
<< metal1 >>
rect -28 15 -18 21
rect -28 12 -22 15
rect -28 11 15 12
rect -28 8 -16 11
rect -17 7 -16 8
rect -12 7 0 11
rect 4 7 10 11
rect 14 7 15 11
rect -17 6 15 7
rect 25 11 41 12
rect 25 7 26 11
rect 30 7 36 11
rect 40 7 41 11
rect 25 6 41 7
rect 51 11 67 12
rect 51 7 52 11
rect 56 7 62 11
rect 66 7 67 11
rect 51 6 67 7
rect 78 11 94 12
rect 78 7 79 11
rect 83 7 89 11
rect 93 7 94 11
rect 78 6 94 7
rect -25 4 -20 5
rect -25 0 -24 4
rect -25 -3 -20 0
rect -1 -3 15 -2
rect -25 -7 -16 -3
rect -12 -7 -11 -3
rect -25 -8 -11 -7
rect -1 -7 0 -3
rect 4 -7 10 -3
rect 14 -7 15 -3
rect -1 -8 15 -7
rect 25 -3 41 -2
rect 25 -7 26 -3
rect 30 -7 36 -3
rect 40 -7 41 -3
rect 25 -8 41 -7
rect 51 -3 67 -2
rect 51 -7 52 -3
rect 56 -7 62 -3
rect 66 -7 67 -3
rect 51 -8 67 -7
rect 78 -3 94 -2
rect 78 -7 79 -3
rect 83 -7 89 -3
rect 93 -7 94 -3
rect 78 -8 94 -7
rect 9 -12 15 -8
rect 9 -16 10 -12
rect 14 -16 15 -12
rect 35 -12 41 -8
rect 35 -16 36 -12
rect 40 -16 41 -12
rect 61 -12 67 -8
rect 61 -16 62 -12
rect 66 -16 67 -12
rect 88 -11 94 -8
rect 88 -12 111 -11
rect 88 -16 89 -12
rect 93 -16 106 -12
rect 110 -16 111 -12
rect 115 -12 121 -11
rect 115 -16 116 -12
rect 120 -16 121 -12
rect 115 -17 121 -16
rect 9 -26 15 -25
rect 9 -30 10 -26
rect 14 -30 15 -26
rect 9 -33 15 -30
rect 35 -26 41 -25
rect 35 -30 36 -26
rect 40 -30 41 -26
rect 35 -33 41 -30
rect 61 -26 67 -25
rect 61 -30 62 -26
rect 66 -30 67 -26
rect 61 -33 67 -30
rect 88 -26 94 -25
rect 88 -30 89 -26
rect 93 -30 94 -26
rect 88 -33 94 -30
rect 105 -26 123 -25
rect 105 -30 106 -26
rect 110 -30 116 -26
rect 120 -30 123 -26
rect 105 -31 123 -30
<< m2contact >>
rect -18 15 -12 21
rect 115 -11 121 -5
rect 9 -39 15 -33
rect 35 -39 41 -33
rect 61 -39 67 -33
rect 88 -39 94 -33
<< metal2 >>
rect -28 15 -18 21
rect -12 15 123 21
rect 97 -11 115 -5
rect 9 -33 15 -25
rect 35 -33 41 -25
rect 61 -33 67 -25
rect 88 -33 94 -25
rect 97 -33 103 -11
rect 115 -16 121 -11
rect -28 -39 9 -33
rect 15 -39 35 -33
rect 41 -39 61 -33
rect 67 -39 88 -33
rect 94 -39 123 -33
<< labels >>
rlabel polysilicon -28 -1 -26 5 3 Iin
rlabel metal1 121 -31 123 -25 8 Iout
rlabel metal2 -28 -39 -22 -33 2 ground
rlabel metal2 -28 15 -22 21 4 Vdd
<< end >>
