magic
tech scmos
timestamp 1418087466
<< ptransistor >>
rect -19 19 -9 29
rect 7 19 17 29
rect 20 19 30 29
rect 33 19 43 29
rect 46 19 56 29
rect 59 19 69 29
rect 72 19 82 29
rect 86 26 96 29
rect 85 21 96 26
rect 86 19 96 21
rect 99 19 109 29
rect 20 0 30 10
rect 46 0 56 10
rect 72 0 82 10
rect 99 0 109 10
rect 121 0 131 10
rect 135 0 145 10
<< pdiffusion >>
rect -19 36 -9 37
rect -19 30 -17 36
rect -11 30 -9 36
rect -19 29 -9 30
rect 7 36 17 37
rect 7 30 9 36
rect 15 30 17 36
rect 7 29 17 30
rect 20 36 30 37
rect 20 30 22 36
rect 28 30 30 36
rect 20 29 30 30
rect 33 36 43 37
rect 33 30 35 36
rect 41 30 43 36
rect 33 29 43 30
rect 46 36 56 37
rect 46 30 48 36
rect 54 30 56 36
rect 46 29 56 30
rect 59 36 69 37
rect 59 30 61 36
rect 67 30 69 36
rect 59 29 69 30
rect 72 36 82 37
rect 72 30 74 36
rect 80 30 82 36
rect 72 29 82 30
rect 86 36 96 37
rect 86 30 88 36
rect 94 30 96 36
rect 86 29 96 30
rect 99 36 109 37
rect 99 30 101 36
rect 107 30 109 36
rect 99 29 109 30
rect -19 18 -9 19
rect -19 12 -17 18
rect -11 12 -9 18
rect -19 11 -9 12
rect 7 18 17 19
rect 7 12 9 18
rect 15 12 17 18
rect 7 11 17 12
rect 20 18 30 19
rect 20 12 22 18
rect 28 12 30 18
rect 20 10 30 12
rect 33 18 43 19
rect 33 12 35 18
rect 41 12 43 18
rect 33 11 43 12
rect 46 18 56 19
rect 46 12 48 18
rect 54 12 56 18
rect 46 10 56 12
rect 59 18 69 19
rect 59 12 61 18
rect 67 12 69 18
rect 59 11 69 12
rect 72 18 82 19
rect 72 12 74 18
rect 80 12 82 18
rect 72 10 82 12
rect 86 18 96 19
rect 86 12 88 18
rect 94 12 96 18
rect 86 11 96 12
rect 99 18 109 19
rect 99 12 101 18
rect 107 12 109 18
rect 99 10 109 12
rect 121 17 131 18
rect 121 11 123 17
rect 129 11 131 17
rect 121 10 131 11
rect 135 17 145 18
rect 135 11 137 17
rect 143 11 145 17
rect 135 10 145 11
rect 20 -1 30 0
rect 20 -7 22 -1
rect 28 -7 30 -1
rect 20 -8 30 -7
rect 46 -1 56 0
rect 46 -7 48 -1
rect 54 -7 56 -1
rect 46 -8 56 -7
rect 72 -1 82 0
rect 72 -7 74 -1
rect 80 -7 82 -1
rect 72 -8 82 -7
rect 99 -1 109 0
rect 99 -7 101 -1
rect 107 -7 109 -1
rect 99 -8 109 -7
rect 121 -1 131 0
rect 121 -7 123 -1
rect 129 -7 131 -1
rect 121 -8 131 -7
rect 135 -1 145 0
rect 135 -7 137 -1
rect 143 -7 145 -1
rect 135 -8 145 -7
<< pdcontact >>
rect -17 30 -11 36
rect 9 30 15 36
rect 22 30 28 36
rect 35 30 41 36
rect 48 30 54 36
rect 61 30 67 36
rect 74 30 80 36
rect 88 30 94 36
rect 101 30 107 36
rect -17 12 -11 18
rect 9 12 15 18
rect 22 12 28 18
rect 35 12 41 18
rect 48 12 54 18
rect 61 12 67 18
rect 74 12 80 18
rect 88 12 94 18
rect 101 12 107 18
rect 123 11 129 17
rect 137 11 143 17
rect 22 -7 28 -1
rect 48 -7 54 -1
rect 74 -7 80 -1
rect 101 -7 107 -1
rect 123 -7 129 -1
rect 137 -7 143 -1
<< polysilicon >>
rect -29 27 -19 29
rect -29 21 -27 27
rect -21 21 -19 27
rect -29 19 -19 21
rect -9 19 7 29
rect 17 19 20 29
rect 30 19 33 29
rect 43 19 46 29
rect 56 19 59 29
rect 69 19 72 29
rect 82 26 86 29
rect 82 21 85 26
rect 82 19 86 21
rect 96 19 99 29
rect 109 19 111 29
rect -6 10 4 19
rect -6 0 20 10
rect 30 0 46 10
rect 56 0 72 10
rect 82 0 99 10
rect 109 0 121 10
rect 131 0 135 10
rect 145 0 147 10
<< polycontact >>
rect -27 21 -21 27
<< metal1 >>
rect -30 39 -17 45
rect -29 36 -22 39
rect -29 30 -17 36
rect -11 30 9 36
rect 15 30 22 36
rect 28 30 30 36
rect 33 30 35 36
rect 41 30 48 36
rect 54 30 56 36
rect 59 30 61 36
rect 67 30 74 36
rect 80 30 82 36
rect 86 30 88 36
rect 94 30 101 36
rect 107 30 109 36
rect 35 26 41 30
rect 61 26 67 30
rect 88 26 94 30
rect -27 18 -21 21
rect 22 21 41 26
rect 48 21 67 26
rect 74 21 94 26
rect 22 18 28 21
rect 48 18 54 21
rect 74 18 80 21
rect -27 12 -17 18
rect 15 12 22 18
rect 41 12 48 18
rect 67 12 74 18
rect 94 12 101 18
rect 137 17 143 19
rect 107 12 123 17
rect 105 11 123 12
rect 14 -7 22 -1
rect 28 -7 48 -1
rect 54 -7 74 -1
rect 80 -7 101 -1
rect 129 -7 137 -1
<< m2contact >>
rect -17 39 -11 45
rect 137 19 143 26
rect 8 -7 14 -1
<< metal2 >>
rect -31 39 -17 45
rect -11 39 149 45
rect -17 30 -11 39
rect 9 30 15 36
rect 22 30 28 36
rect 35 30 41 36
rect 48 30 54 36
rect 61 30 67 36
rect 74 30 80 36
rect 88 30 94 36
rect 101 30 107 36
rect 113 19 137 26
rect 143 19 149 26
rect 113 -1 119 19
rect 137 11 143 19
rect -31 -7 8 -1
rect 14 -7 119 -1
<< labels >>
rlabel metal2 146 20 148 24 7 Gnd
rlabel metal2 146 40 148 44 6 Vdd
rlabel metal2 -29 -6 -27 -2 2 Gnd
<< end >>
