magic
tech scmos
timestamp 1417635104
<< ntransistor >>
rect 3 0 9 6
rect 15 0 21 6
rect 35 0 41 6
rect 47 0 53 6
rect 67 0 73 6
rect 79 0 85 6
rect 99 5 105 11
rect 99 -19 105 -13
<< ptransistor >>
rect 3 55 9 61
rect 15 55 21 61
rect 35 55 41 61
rect 47 55 53 61
rect 67 55 73 61
rect 79 55 85 61
rect 99 55 105 61
rect 111 55 117 61
rect 131 55 137 61
rect 143 55 149 61
<< ndiffusion >>
rect 94 10 99 11
rect 98 6 99 10
rect -2 5 3 6
rect 2 1 3 5
rect -2 0 3 1
rect 9 5 15 6
rect 9 1 10 5
rect 14 1 15 5
rect 9 0 15 1
rect 21 5 26 6
rect 21 1 22 5
rect 21 0 26 1
rect 30 5 35 6
rect 34 1 35 5
rect 30 0 35 1
rect 41 5 47 6
rect 41 1 42 5
rect 46 1 47 5
rect 41 0 47 1
rect 53 5 58 6
rect 53 1 54 5
rect 53 0 58 1
rect 62 5 67 6
rect 66 1 67 5
rect 62 0 67 1
rect 73 5 79 6
rect 73 1 74 5
rect 78 1 79 5
rect 73 0 79 1
rect 85 5 90 6
rect 94 5 99 6
rect 105 10 110 11
rect 105 6 106 10
rect 105 5 110 6
rect 85 1 86 5
rect 85 0 90 1
rect 94 -14 99 -13
rect 98 -18 99 -14
rect 94 -19 99 -18
rect 105 -14 110 -13
rect 105 -18 106 -14
rect 105 -19 110 -18
<< pdiffusion >>
rect 42 83 46 87
rect 62 83 66 87
rect 86 83 90 87
rect 126 83 130 87
rect 150 83 154 87
rect 10 61 14 65
rect -2 60 3 61
rect 2 56 3 60
rect -2 55 3 56
rect 9 60 15 61
rect 9 56 10 60
rect 14 56 15 60
rect 9 55 15 56
rect 21 60 26 61
rect 21 56 22 60
rect 21 55 26 56
rect 30 60 35 61
rect 34 56 35 60
rect 30 55 35 56
rect 41 60 47 61
rect 41 56 42 60
rect 46 56 47 60
rect 41 55 47 56
rect 53 60 58 61
rect 53 56 54 60
rect 53 55 58 56
rect 62 60 67 61
rect 66 56 67 60
rect 62 55 67 56
rect 73 60 79 61
rect 73 56 74 60
rect 78 56 79 60
rect 73 55 79 56
rect 85 60 90 61
rect 85 56 86 60
rect 85 55 90 56
rect 94 60 99 61
rect 98 56 99 60
rect 94 55 99 56
rect 105 60 111 61
rect 105 56 106 60
rect 110 56 111 60
rect 105 55 111 56
rect 117 60 122 61
rect 117 56 118 60
rect 117 55 122 56
rect 126 60 131 61
rect 130 56 131 60
rect 126 55 131 56
rect 137 60 143 61
rect 137 56 138 60
rect 142 56 143 60
rect 137 55 143 56
rect 149 60 154 61
rect 149 56 150 60
rect 149 55 154 56
<< ndcontact >>
rect 94 6 98 10
rect -2 1 2 5
rect 10 1 14 5
rect 22 1 26 5
rect 30 1 34 5
rect 42 1 46 5
rect 54 1 58 5
rect 62 1 66 5
rect 74 1 78 5
rect 106 6 110 10
rect 86 1 90 5
rect 94 -18 98 -14
rect 106 -18 110 -14
<< pdcontact >>
rect -2 56 2 60
rect 10 56 14 60
rect 22 56 26 60
rect 30 56 34 60
rect 42 56 46 60
rect 54 56 58 60
rect 62 56 66 60
rect 74 56 78 60
rect 86 56 90 60
rect 94 56 98 60
rect 106 56 110 60
rect 118 56 122 60
rect 126 56 130 60
rect 138 56 142 60
rect 150 56 154 60
<< psubstratepcontact >>
rect 1 -28 39 -24
rect 49 -28 71 -24
rect 82 -28 115 -24
rect 126 -28 153 -24
<< nsubstratencontact >>
rect 0 83 6 87
rect 17 83 38 87
rect 50 83 58 87
rect 70 83 82 87
rect 94 83 121 87
rect 134 83 146 87
<< polysilicon >>
rect 3 61 9 63
rect 15 61 21 63
rect 35 61 41 63
rect 47 61 53 63
rect 67 61 73 63
rect 79 61 85 63
rect 99 61 105 63
rect 111 61 117 63
rect 131 61 137 63
rect 143 61 149 63
rect 3 53 9 55
rect 3 49 4 53
rect 8 52 9 53
rect 15 52 21 55
rect 8 49 21 52
rect 35 54 41 55
rect 39 53 41 54
rect 47 53 53 55
rect 67 53 73 55
rect 39 50 73 53
rect 35 49 73 50
rect 79 53 85 55
rect 99 53 105 55
rect 111 53 117 55
rect 83 49 85 53
rect 115 49 117 53
rect 131 53 137 55
rect 135 49 137 53
rect 143 53 149 55
rect 143 49 146 53
rect 99 11 105 13
rect 3 6 9 8
rect 15 6 21 8
rect 35 6 41 8
rect 47 6 53 8
rect 67 6 73 8
rect 79 6 85 8
rect 3 -2 9 0
rect 3 -3 4 -2
rect 8 -3 9 -2
rect 15 -2 21 0
rect 15 -3 16 -2
rect 20 -3 21 -2
rect 35 -2 41 0
rect 47 -2 53 0
rect 39 -3 41 -2
rect 67 -2 73 0
rect 79 -2 85 0
rect 99 -2 105 5
rect 71 -6 83 -2
rect 99 -6 100 -2
rect 104 -6 105 -2
rect 99 -13 105 -6
rect 99 -21 105 -19
<< polycontact >>
rect 99 63 103 67
rect 113 63 117 67
rect 4 49 8 53
rect 35 50 39 54
rect 79 49 83 53
rect 111 49 115 53
rect 131 49 135 53
rect 146 49 150 53
rect 4 -6 8 -2
rect 16 -6 20 -2
rect 35 -6 39 -2
rect 49 -6 53 -2
rect 67 -6 71 -2
rect 83 -6 87 -2
rect 100 -6 104 -2
<< metal1 >>
rect -3 87 156 88
rect -3 83 0 87
rect 6 83 10 87
rect 14 83 17 87
rect 38 83 42 87
rect 46 83 50 87
rect 58 83 62 87
rect 66 83 70 87
rect 82 83 86 87
rect 90 83 94 87
rect 121 83 126 87
rect 130 83 134 87
rect 146 83 150 87
rect 154 83 156 87
rect -3 82 156 83
rect 78 75 106 79
rect -3 68 103 72
rect 99 67 103 68
rect 10 60 14 61
rect 42 60 46 61
rect 62 60 66 61
rect -2 53 2 56
rect 2 49 4 53
rect 22 39 26 56
rect 74 60 78 61
rect 113 68 142 72
rect 113 67 117 68
rect 86 60 90 61
rect 106 60 110 61
rect 126 60 130 61
rect 122 56 123 60
rect 138 60 142 68
rect 150 60 154 61
rect 30 55 34 56
rect 54 55 58 56
rect 34 51 35 54
rect 30 50 35 51
rect 94 53 98 56
rect 119 55 123 56
rect 78 49 79 53
rect 111 46 115 49
rect 131 39 135 49
rect 22 35 54 39
rect 58 35 135 39
rect 145 49 146 53
rect 141 32 145 49
rect 2 28 79 32
rect 83 28 145 32
rect 58 21 156 25
rect 10 13 34 17
rect 66 14 156 18
rect -2 5 2 6
rect 10 5 14 13
rect 22 5 26 6
rect 30 5 34 13
rect 54 5 58 6
rect 62 5 66 6
rect 86 5 90 6
rect 42 0 46 1
rect -3 -6 4 -2
rect 16 -9 20 -6
rect -3 -13 20 -9
rect 74 0 78 1
rect 53 -6 67 -2
rect 94 5 98 6
rect 106 5 110 6
rect 86 -2 90 1
rect 87 -6 100 -2
rect 35 -16 39 -6
rect -3 -20 39 -16
rect 94 -14 98 -13
rect 106 -14 110 -13
rect 94 -23 98 -18
rect -3 -24 156 -23
rect -3 -28 1 -24
rect 39 -28 42 -24
rect 46 -28 49 -24
rect 71 -28 74 -24
rect 78 -28 82 -24
rect 115 -28 119 -24
rect 123 -28 126 -24
rect 153 -28 156 -24
rect -3 -29 156 -28
<< m2contact >>
rect 10 83 14 87
rect 42 83 46 87
rect 62 83 66 87
rect 86 83 90 87
rect 126 83 130 87
rect 150 83 154 87
rect 74 75 78 79
rect 106 75 110 79
rect 10 61 14 65
rect 42 61 46 65
rect 62 61 66 65
rect -2 49 2 53
rect 74 61 78 65
rect 86 61 90 65
rect 106 61 110 65
rect 126 61 130 65
rect 150 61 154 65
rect 30 51 34 55
rect 54 51 58 55
rect 74 49 78 53
rect 94 49 98 53
rect 119 51 123 55
rect 111 42 115 46
rect 54 35 58 39
rect 141 49 145 53
rect -2 28 2 32
rect 79 28 83 32
rect 54 21 58 25
rect 62 14 66 18
rect -2 6 2 10
rect 22 6 26 10
rect 54 6 58 10
rect 62 6 66 10
rect 86 6 90 10
rect 42 -4 46 0
rect 74 -4 78 0
rect 94 1 98 5
rect 106 1 110 5
rect 94 -13 98 -9
rect 106 -13 110 -9
rect 42 -28 46 -24
rect 74 -28 78 -24
rect 119 -28 123 -24
<< metal2 >>
rect 10 65 14 83
rect 42 65 46 83
rect 42 60 46 61
rect 62 65 66 83
rect 74 65 78 75
rect 86 65 90 83
rect 106 65 110 75
rect 126 65 130 83
rect 150 65 154 83
rect 62 60 66 61
rect 86 60 90 61
rect -2 32 2 49
rect -2 10 2 28
rect 22 51 30 55
rect 58 51 66 55
rect 22 10 26 51
rect 54 25 58 35
rect 54 10 58 21
rect 62 18 66 51
rect 74 40 78 49
rect 86 49 94 53
rect 74 36 83 40
rect 79 32 83 36
rect 62 10 66 14
rect 86 10 90 49
rect 111 5 115 42
rect 42 -24 46 -4
rect 74 -24 78 -4
rect 94 -9 98 1
rect 110 1 115 5
rect 106 -9 110 1
rect 119 -24 123 51
<< labels >>
rlabel metal1 -3 69 -2 71 3 Vcm
rlabel metal1 19 -29 23 -28 1 GND
rlabel metal1 -3 -5 -2 -3 3 V1
rlabel metal1 -3 -12 -2 -10 3 V2
rlabel metal1 -3 -19 -2 -17 3 Vb
rlabel metal1 155 22 156 24 7 Vout+
rlabel metal1 155 15 156 17 7 Vout-
<< end >>
