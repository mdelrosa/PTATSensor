magic
tech scmos
timestamp 1418681314
<< ntransistor >>
rect -6 -105 394 -101
rect 399 -105 800 -101
rect 804 -105 844 -101
rect -45 -513 -41 -113
rect -1 -513 3 -113
rect 311 -244 324 -234
<< ptransistor >>
rect 108 -46 138 -36
rect 156 -46 166 -36
rect 175 -46 185 -36
rect 191 -46 204 -36
<< ndiffusion >>
rect 836 -95 844 -94
rect -6 -96 394 -95
rect -6 -100 -5 -96
rect 393 -100 394 -96
rect -6 -101 394 -100
rect 399 -96 800 -95
rect 399 -100 400 -96
rect 798 -100 800 -96
rect 399 -101 800 -100
rect 804 -96 844 -95
rect 804 -100 811 -96
rect 837 -100 844 -96
rect 804 -101 844 -100
rect -49 -102 -37 -101
rect -49 -110 -48 -102
rect -38 -110 -37 -102
rect -49 -111 -37 -110
rect -45 -113 -41 -111
rect -6 -106 394 -105
rect -6 -110 -5 -106
rect 393 -110 394 -106
rect -6 -111 394 -110
rect 399 -106 800 -105
rect 399 -110 400 -106
rect 798 -110 800 -106
rect 399 -111 800 -110
rect 804 -106 844 -105
rect 804 -110 811 -106
rect 837 -110 844 -106
rect 804 -111 844 -110
rect -1 -113 3 -111
rect 404 -112 408 -111
rect 311 -224 324 -223
rect 311 -233 312 -224
rect 323 -233 324 -224
rect 311 -234 324 -233
rect 311 -245 324 -244
rect 311 -254 312 -245
rect 323 -254 324 -245
rect 311 -255 324 -254
rect -45 -515 -41 -513
rect -1 -514 3 -513
rect -5 -515 7 -514
rect -49 -516 -37 -515
rect -49 -520 -48 -516
rect -38 -520 -37 -516
rect -5 -519 -4 -515
rect 6 -519 7 -515
rect -5 -520 7 -519
rect -49 -521 -37 -520
<< pdiffusion >>
rect 156 -30 166 -29
rect 108 -31 138 -30
rect 108 -35 109 -31
rect 137 -35 138 -31
rect 108 -36 138 -35
rect 156 -35 157 -30
rect 165 -35 166 -30
rect 156 -36 166 -35
rect 175 -30 185 -29
rect 175 -35 176 -30
rect 184 -35 185 -30
rect 175 -36 185 -35
rect 191 -30 204 -29
rect 191 -35 192 -30
rect 203 -35 204 -30
rect 191 -36 204 -35
rect 108 -47 138 -46
rect 108 -51 109 -47
rect 137 -51 138 -47
rect 108 -52 138 -51
rect 156 -48 166 -46
rect 156 -53 157 -48
rect 165 -53 166 -48
rect 156 -54 166 -53
rect 175 -48 185 -46
rect 175 -53 176 -48
rect 184 -53 185 -48
rect 175 -54 185 -53
rect 191 -48 204 -46
rect 191 -53 192 -48
rect 203 -53 204 -48
rect 191 -54 204 -53
<< ndcontact >>
rect -5 -100 393 -96
rect 400 -100 798 -96
rect 811 -100 837 -96
rect -48 -110 -38 -102
rect -5 -110 393 -106
rect 400 -110 798 -106
rect 811 -110 837 -106
rect 312 -233 323 -224
rect 312 -254 323 -245
rect -48 -520 -38 -516
rect -4 -519 6 -515
<< pdcontact >>
rect 109 -35 137 -31
rect 157 -35 165 -30
rect 176 -35 184 -30
rect 192 -35 203 -30
rect 109 -51 137 -47
rect 157 -53 165 -48
rect 176 -53 184 -48
rect 192 -53 203 -48
<< polysilicon >>
rect 105 -46 108 -36
rect 138 -46 156 -36
rect 166 -46 175 -36
rect 185 -46 191 -36
rect 204 -46 210 -36
rect 143 -48 151 -46
rect 143 -53 144 -48
rect 150 -53 151 -48
rect 143 -54 151 -53
rect -36 -103 -27 -102
rect -36 -109 -35 -103
rect -28 -109 -27 -103
rect -9 -105 -6 -101
rect 394 -105 399 -101
rect 800 -105 804 -101
rect 844 -105 847 -101
rect -36 -113 -27 -109
rect -49 -513 -45 -113
rect -41 -513 -1 -113
rect 3 -234 7 -113
rect 3 -244 311 -234
rect 324 -244 327 -234
rect 3 -513 7 -244
<< polycontact >>
rect 144 -53 150 -48
rect -35 -109 -28 -103
<< metal1 >>
rect 100 -31 157 -30
rect 100 -35 109 -31
rect 137 -35 157 -31
rect 165 -35 176 -30
rect 184 -35 192 -30
rect 203 -35 213 -30
rect -49 -51 109 -48
rect 176 -48 184 -47
rect 137 -51 138 -48
rect -49 -52 138 -51
rect -49 -102 -38 -52
rect 143 -53 144 -48
rect 150 -53 157 -48
rect 165 -53 166 -48
rect 156 -92 166 -53
rect 176 -61 184 -53
rect 191 -53 192 -48
rect 203 -53 857 -48
rect 191 -55 857 -53
rect 191 -56 454 -55
rect 176 -64 833 -61
rect 175 -67 833 -64
rect -5 -96 798 -92
rect 393 -100 400 -96
rect 811 -94 833 -67
rect 811 -95 837 -94
rect 811 -96 839 -95
rect 837 -100 839 -96
rect -5 -101 798 -100
rect -50 -110 -48 -102
rect -38 -103 -27 -102
rect -38 -109 -35 -103
rect -28 -109 -27 -103
rect 386 -106 409 -105
rect -38 -110 -27 -109
rect 393 -110 400 -106
rect -50 -111 -27 -110
rect 386 -111 409 -110
rect 811 -116 831 -110
rect 312 -224 856 -223
rect 323 -233 856 -224
rect 312 -257 323 -254
rect 312 -263 320 -257
rect 313 -511 320 -263
rect 313 -515 321 -511
rect 347 -515 372 -511
rect -49 -516 -29 -515
rect -49 -520 -48 -516
rect -38 -520 -29 -516
rect -18 -519 -4 -515
rect 6 -519 266 -515
rect -18 -520 266 -519
rect 277 -520 372 -515
rect 313 -521 321 -520
rect 347 -523 372 -520
<< m2contact >>
rect 93 -35 100 -30
rect 213 -35 220 -30
rect 811 -125 832 -116
rect -29 -523 -18 -515
rect 266 -523 277 -515
<< metal2 >>
rect -59 -30 857 -27
rect -59 -35 93 -30
rect 100 -35 213 -30
rect 220 -35 857 -30
rect -59 -36 857 -35
rect 811 -116 832 -106
rect 811 -512 832 -125
rect 442 -514 867 -512
rect -50 -515 867 -514
rect -50 -523 -29 -515
rect -18 -523 266 -515
rect 277 -523 867 -515
rect -50 -524 867 -523
rect 442 -525 867 -524
rect 471 -526 488 -525
<< labels >>
rlabel metal2 852 -35 855 -29 6 Vdd
rlabel metal1 852 -54 855 -48 7 I_push
rlabel metal1 851 -231 855 -224 7 I_pull
rlabel metal2 860 -523 865 -515 7 Gnd
<< end >>
