magic
tech scmos
timestamp 1417640631
<< nwell >>
rect -77 -94 -39 -56
<< ntransistor >>
rect -27 9 -21 15
rect -7 9 -1 15
rect -27 -36 -21 -30
rect -7 -36 -1 -30
<< ndiffusion >>
rect -27 21 -21 22
rect -27 17 -26 21
rect -22 17 -21 21
rect -27 15 -21 17
rect -7 21 -1 22
rect -7 17 -6 21
rect -2 17 -1 21
rect -7 15 -1 17
rect -27 7 -21 9
rect -27 3 -26 7
rect -22 3 -21 7
rect -27 2 -21 3
rect -7 7 -1 9
rect -7 3 -6 7
rect -2 3 -1 7
rect -7 2 -1 3
rect -27 -24 -21 -23
rect -27 -28 -26 -24
rect -22 -28 -21 -24
rect -27 -30 -21 -28
rect -7 -24 -1 -23
rect -7 -28 -6 -24
rect -2 -28 -1 -24
rect -7 -30 -1 -28
rect -27 -38 -21 -36
rect -27 -42 -26 -38
rect -22 -42 -21 -38
rect -27 -43 -21 -42
rect -7 -38 -1 -36
rect -7 -42 -6 -38
rect -2 -42 -1 -38
rect -7 -43 -1 -42
<< pdiffusion >>
rect -64 -70 -52 -69
rect -64 -80 -63 -70
rect -53 -80 -52 -70
rect -64 -81 -52 -80
<< ndcontact >>
rect -26 17 -22 21
rect -6 17 -2 21
rect -26 3 -22 7
rect -6 3 -2 7
rect -26 -28 -22 -24
rect -6 -28 -2 -24
rect -26 -42 -22 -38
rect -6 -42 -2 -38
<< pdcontact >>
rect -63 -80 -53 -70
<< psubstratepdiff >>
rect -86 -48 -30 -47
rect -86 -52 -85 -48
rect -31 -52 -30 -48
rect -86 -53 -30 -52
rect -86 -55 -80 -53
rect -86 -95 -85 -55
rect -81 -95 -80 -55
rect -36 -55 -30 -53
rect -36 -67 -35 -55
rect -31 -67 -30 -55
rect -36 -84 -30 -67
rect -86 -97 -80 -95
rect -36 -95 -35 -84
rect -31 -95 -30 -84
rect -36 -97 -30 -95
rect -86 -98 -30 -97
rect -86 -102 -85 -98
rect -31 -102 -30 -98
rect -86 -103 -30 -102
<< nsubstratendiff >>
rect -74 -60 -42 -59
rect -74 -64 -73 -60
rect -43 -64 -42 -60
rect -74 -65 -42 -64
rect -74 -67 -68 -65
rect -74 -83 -73 -67
rect -69 -83 -68 -67
rect -48 -77 -42 -65
rect -74 -85 -68 -83
rect -48 -83 -47 -77
rect -43 -83 -42 -77
rect -48 -85 -42 -83
rect -74 -86 -42 -85
rect -74 -90 -73 -86
rect -43 -90 -42 -86
rect -74 -91 -42 -90
<< psubstratepcontact >>
rect -85 -52 -31 -48
rect -85 -95 -81 -55
rect -35 -67 -31 -55
rect -35 -95 -31 -84
rect -85 -102 -31 -98
<< nsubstratencontact >>
rect -73 -64 -43 -60
rect -73 -83 -69 -67
rect -47 -83 -43 -77
rect -73 -90 -43 -86
<< polysilicon >>
rect -85 9 -27 15
rect -21 9 -7 15
rect -1 9 46 15
rect -85 -36 -27 -30
rect -21 -36 -7 -30
rect -1 -36 46 -30
<< metal1 >>
rect -7 32 8 38
rect -36 23 -21 29
rect -44 -38 -39 -15
rect -36 -23 -30 23
rect -27 21 -21 23
rect -27 17 -26 21
rect -22 17 -21 21
rect -7 21 -1 32
rect -7 17 -6 21
rect -2 17 -1 21
rect -27 3 -26 7
rect -22 3 -13 7
rect -27 0 -13 3
rect -36 -24 -21 -23
rect -36 -28 -26 -24
rect -22 -28 -21 -24
rect -18 -38 -13 0
rect -7 3 -6 7
rect -2 3 -1 7
rect -7 -9 -1 3
rect 2 -23 8 32
rect -7 -24 8 -23
rect -7 -28 -6 -24
rect -2 -28 8 -24
rect -85 -42 -26 -38
rect -22 -42 -21 -38
rect -85 -43 -21 -42
rect -18 -42 -6 -38
rect -2 -42 46 -38
rect -18 -43 46 -42
rect -85 -55 -81 -52
rect -35 -55 -31 -52
rect -73 -67 -69 -64
rect -27 -70 -21 -43
rect -53 -74 -21 -70
rect -7 -70 -1 -43
rect -7 -74 5 -70
rect -73 -86 -69 -83
rect -43 -81 -23 -77
rect -47 -86 -43 -83
rect -28 -84 -23 -81
rect -85 -98 -81 -95
rect -31 -88 -23 -84
rect -35 -98 -31 -95
rect -28 -107 -23 -88
rect -3 -107 2 -77
rect -28 -112 -16 -107
rect -11 -112 4 -107
<< m2contact >>
rect -13 32 -7 38
rect -21 23 -15 29
rect -44 -15 -39 -9
rect -7 -15 -1 -9
rect -16 -112 -11 -107
<< metal2 >>
rect -85 32 -13 38
rect -7 32 45 38
rect -85 23 -21 29
rect -15 23 45 29
rect -45 -15 -44 -9
rect -39 -15 -7 -9
rect -86 -112 -16 -107
rect -11 -112 45 -107
use CVBT  CVBT_0
timestamp 1415294909
transform -1 0 61 0 -1 -47
box 0 0 59 56
<< labels >>
rlabel metal1 -28 -73 -27 -71 3 E
rlabel metal1 -28 -80 -27 -78 3 B
rlabel metal1 -28 -87 -27 -85 3 C
rlabel metal1 -85 -43 -83 -38 3 dVbe+
rlabel metal1 44 -43 46 -38 1 dVbe-
rlabel metal2 -84 33 -82 37 4 NI_Iin
rlabel metal2 -84 24 -82 28 3 Iin
rlabel polysilicon -84 10 -82 14 3 clk
rlabel polysilicon -84 -35 -82 -31 3 nclk
rlabel metal2 -85 -111 -83 -107 2 gnd
<< end >>
