magic
tech scmos
timestamp 1418250215
<< ntransistor >>
rect -647 -9 -527 -3
rect -515 -9 -395 -3
rect -379 -9 -259 -3
rect -247 -9 -127 -3
rect -114 -9 6 -3
rect 18 -9 138 -3
rect 151 -9 271 -3
rect 283 -9 403 -3
<< ptransistor >>
rect -647 55 -527 61
rect -515 55 -395 61
rect -379 55 -259 61
rect -247 55 -127 61
rect -114 55 6 61
rect 18 55 138 61
rect 151 55 271 61
rect 284 55 404 61
rect 417 55 537 61
rect 556 55 676 61
<< ndiffusion >>
rect -647 0 -640 1
rect -647 -3 -527 0
rect -515 -1 -402 0
rect -515 -3 -395 -1
rect -372 -1 -259 0
rect -379 -3 -259 -1
rect -240 -1 -127 0
rect -247 -3 -127 -1
rect -107 -1 6 0
rect -114 -3 6 -1
rect 18 -1 132 0
rect 266 0 290 6
rect 18 -3 138 -1
rect 151 -1 396 0
rect 151 -3 271 -1
rect 283 -3 403 -1
rect -647 -11 -527 -9
rect -515 -11 -395 -9
rect -647 -12 -402 -11
rect -531 -17 -510 -12
rect -379 -11 -259 -9
rect -247 -11 -127 -9
rect -379 -12 -127 -11
rect -114 -11 6 -9
rect 18 -11 138 -9
rect -114 -12 138 -11
rect 151 -11 271 -9
rect 283 -11 403 -9
rect 151 -12 403 -11
rect -266 -17 -256 -12
rect -250 -17 -242 -12
rect 1 -15 9 -12
rect 14 -15 23 -12
rect 266 -17 274 -12
rect 280 -17 288 -12
<< pdiffusion >>
rect -531 64 -524 69
rect -647 63 -524 64
rect -518 64 -510 69
rect -265 64 -256 69
rect -518 63 -395 64
rect -647 61 -527 63
rect -515 61 -395 63
rect -379 63 -256 64
rect -250 64 -241 69
rect 1 64 18 68
rect -250 63 -127 64
rect -379 61 -259 63
rect -247 61 -127 63
rect -114 63 18 64
rect 25 63 138 64
rect -114 61 6 63
rect 18 61 138 63
rect 151 63 165 64
rect 267 64 289 69
rect 533 64 543 72
rect 551 64 561 72
rect 172 63 404 64
rect -647 53 -527 55
rect -640 52 -527 53
rect -515 53 -395 55
rect 151 61 271 63
rect 284 61 404 63
rect 417 63 676 64
rect 417 61 537 63
rect 556 61 676 63
rect -379 53 -259 55
rect -515 52 -401 53
rect -372 52 -259 53
rect -247 53 -127 55
rect -247 52 -151 53
rect -144 52 -127 53
rect -114 53 6 55
rect 18 53 138 55
rect -114 52 10 53
rect 1 48 10 52
rect 15 52 138 53
rect 151 53 271 55
rect 15 48 23 52
rect 159 52 271 53
rect 284 53 404 55
rect 284 52 346 53
rect 353 52 404 53
rect 417 53 537 55
rect 556 53 676 55
rect 424 52 676 53
rect 533 45 561 52
<< ndcontact >>
rect -647 1 -640 8
rect -402 -1 -395 6
rect -379 -1 -372 6
rect -247 -1 -240 6
rect -114 -1 -107 6
rect 132 -1 138 5
rect 396 -1 403 6
rect -402 -18 -395 -11
rect -256 -18 -250 -12
rect 9 -17 14 -12
rect 274 -18 280 -12
<< pdcontact >>
rect -524 63 -518 69
rect -256 63 -250 69
rect 18 63 25 70
rect 165 63 172 70
rect 543 64 551 72
rect -647 46 -640 53
rect -401 46 -394 53
rect -379 46 -372 53
rect -151 46 -144 53
rect 10 48 15 53
rect 151 45 159 53
rect 346 46 353 53
rect 417 46 424 53
<< psubstratepcontact >>
rect -660 -49 688 -44
<< nsubstratencontact >>
rect -660 87 688 92
<< polysilicon >>
rect -649 55 -647 61
rect -527 55 -515 61
rect -395 55 -392 61
rect -381 55 -379 61
rect -259 55 -247 61
rect -127 55 -114 61
rect 6 55 9 61
rect 15 55 18 61
rect 138 56 139 61
rect 138 55 145 56
rect 149 55 151 61
rect 271 56 272 61
rect 271 55 278 56
rect 282 55 284 61
rect 404 55 405 61
rect 415 55 417 61
rect 537 55 538 61
rect 554 55 556 61
rect 676 55 678 61
rect -649 -9 -647 -3
rect -527 -9 -525 -3
rect -521 -4 -515 -3
rect -516 -9 -515 -4
rect -395 -9 -392 -3
rect -382 -9 -379 -3
rect -259 -9 -257 -3
rect -253 -9 -247 -3
rect -127 -9 -114 -3
rect 6 -9 18 -3
rect 138 -9 140 -3
rect 147 -9 151 -3
rect 271 -9 283 -3
rect 403 -9 407 -3
<< polycontact >>
rect -656 54 -649 61
rect -388 54 -381 61
rect 139 56 145 62
rect 272 56 278 62
rect 405 55 411 61
rect 538 55 544 61
rect 678 55 685 62
rect -655 -9 -649 -3
rect -521 -9 -516 -4
rect -388 -9 -382 -3
rect 140 -9 147 -2
<< metal1 >>
rect -661 92 689 93
rect -661 87 -660 92
rect 688 87 689 92
rect -661 86 689 87
rect -661 75 -655 81
rect -524 69 -518 86
rect -256 69 -250 86
rect -656 47 -647 54
rect -388 53 -381 54
rect 10 53 15 86
rect 25 63 27 70
rect 163 63 165 70
rect 272 62 278 75
rect 543 72 551 86
rect -647 35 -640 46
rect -388 47 -379 53
rect -401 45 -394 46
rect -647 8 -640 28
rect -379 25 -372 46
rect 123 56 139 62
rect -402 6 -395 18
rect -247 6 -240 38
rect -151 15 -144 46
rect 123 35 130 56
rect 405 53 411 55
rect 140 45 151 53
rect 405 46 417 53
rect -114 6 -107 8
rect 140 5 147 45
rect 138 -1 147 5
rect -661 -9 -655 -3
rect -521 -19 -516 -9
rect -661 -25 -655 -19
rect -402 -19 -395 -18
rect -388 -31 -382 -9
rect -379 -19 -372 -1
rect 140 -2 147 -1
rect -661 -37 -655 -31
rect -256 -43 -250 -18
rect 9 -43 14 -17
rect 274 -43 280 -18
rect 346 -43 353 46
rect 417 6 424 46
rect 538 25 544 55
rect 662 55 678 61
rect 662 35 669 55
rect 681 38 688 45
rect 681 8 688 15
rect 403 -1 424 6
rect -661 -44 689 -43
rect -661 -49 -660 -44
rect 688 -49 689 -44
rect -661 -50 689 -49
<< m2contact >>
rect -655 75 -649 81
rect 272 75 278 81
rect 27 63 34 70
rect 156 63 163 70
rect -401 38 -394 45
rect -647 28 -640 35
rect -402 18 -395 25
rect -379 18 -372 25
rect -247 38 -240 45
rect 123 28 130 35
rect -151 8 -144 15
rect -114 8 -107 15
rect -655 -25 -649 -19
rect -522 -25 -516 -19
rect -402 -26 -395 -19
rect -379 -26 -372 -19
rect -655 -37 -649 -31
rect -388 -37 -382 -31
rect 674 38 681 45
rect 662 28 669 35
rect 537 18 544 25
rect 674 8 681 15
<< metal2 >>
rect -649 75 272 81
rect 34 63 156 70
rect -394 38 -247 45
rect -240 38 674 45
rect -640 28 123 35
rect 130 28 662 35
rect -395 18 -379 25
rect -372 18 537 25
rect -144 8 -114 15
rect -107 8 674 15
rect -649 -25 -522 -19
rect -395 -26 -379 -19
rect -649 -37 -388 -31
<< labels >>
rlabel metal1 681 38 688 45 7 Vout+
rlabel metal1 681 8 688 15 7 Vout-
rlabel metal1 -661 75 -655 81 3 Vcm
rlabel metal1 -661 -9 -655 -3 3 V1
rlabel metal1 -661 -25 -655 -19 3 V2
rlabel metal1 -661 -37 -655 -31 3 Vb
rlabel metal1 -661 86 689 93 5 VDD
rlabel metal1 -661 -50 689 -43 1 GND
<< end >>
